0
0 1 0 1 0 g 1 c
0 2 4 0 0 g c
0 2 2 1 0 g c
7 0 5 0 0 g c
4 5 0 3 0 10 0 4 2 8 1 9 0 6 3 11 2 12 3 3 5 7 3 10 4 2 1 9 2 5 2 6 4 11 1 8 1 4
0
